`include "header.v"

module alu(
    
);

endmodule