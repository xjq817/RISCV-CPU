`include "header.v"

module LSB(
    input  wire  clk,
    input  wire  rst,
    input  wire  rdy,
    input  wire  jump_wrong,
//MemoryController
//decoder
//RS
//ROB
//for all
);


endmodule