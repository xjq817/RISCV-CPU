`include "header.v"

module LSB(
    
);

endmodule