`include "header.v"

module IF(
    
);

endmodule