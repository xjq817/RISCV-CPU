`include "header.v"

module ROB(
    
);

endmodule