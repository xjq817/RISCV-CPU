`include "header.v"

module RS(
    
);

endmodule