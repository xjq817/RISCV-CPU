`include "header.v"

module MemoryController (
    
);



endmodule