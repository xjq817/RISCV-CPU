`include "define.v"

module decoder(
    input  wire  clk,
    input  wire  rst,
    input  wire  rdy,
);

    
endmodule